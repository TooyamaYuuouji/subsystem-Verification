`define TIMER0_OFFSET 16'h0000
`define TIMER0_CTRL_OFFSET `TIMER0_OFFSET+16'h0000
`define TIMER0_VALUE_OFFSET 16'h0004
`define TIMER0_RELOAD_OFFSET 16'h0008
`define TIMER0_INTCLEAR_OFFSET 16'h000C

`define APB_TEST_SLAVE_OFFSET 16'hB000
`define APB_TEST_SLAVE_DATA0_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0000
`define APB_TEST_SLAVE_DATA1_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0004
`define APB_TEST_SLAVE_DATA2_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0008
`define APB_TEST_SLAVE_DATA3_OFFSET `APB_TEST_SLAVE_OFFSET+16'h000C