
package top_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "base_test.sv"

endpackage: top_pkg