`define TIMER0_OFFSET 16'h0000
`define TIMER0_CTRL_OFFSET `TIMER0_OFFSET+16'h0000
`define TIMER0_VALUE_OFFSET `TIMER0_OFFSET+16'h0004
`define TIMER0_RELOAD_OFFSET `TIMER0_OFFSET+16'h0008
`define TIMER0_INTCLEAR_OFFSET `TIMER0_OFFSET+16'h000C

`define TIMER1_OFFSET 16'h1000
`define TIMER1_CTRL_OFFSET `TIMER1_OFFSET+16'h0000
`define TIMER1_VALUE_OFFSET `TIMER1_OFFSET+16'h0004
`define TIMER1_RELOAD_OFFSET `TIMER1_OFFSET+16'h0008
`define TIMER1_INTCLEAR_OFFSET `TIMER1_OFFSET+16'h000C

`define DUALTIMER_OFFSET 16'h2000
`define DUALTIMER_TIMER1LOAD_OFFSET `DUALTIMER_OFFSET+16'h0000
`define DUALTIMER_TIMER1VALUE_OFFSET `DUALTIMER_OFFSET+16'h0004
`define DUALTIMER_TIMER1CONTROL_OFFSET `DUALTIMER_OFFSET+16'h0008
`define DUALTIMER_TIMER1INTCLR_OFFSET `DUALTIMER_OFFSET+16'h000C
`define DUALTIMER_TIMER1RIS_OFFSET `DUALTIMER_OFFSET+16'h0010
`define DUALTIMER_TIMER1MIS_OFFSET `DUALTIMER_OFFSET+16'h0014
`define DUALTIMER_TIMER1BGLOAD_OFFSET `DUALTIMER_OFFSET+16'h0018
`define DUALTIMER_TIMER2LOAD_OFFSET `DUALTIMER_OFFSET+16'h0020
`define DUALTIMER_TIMER2VALUE_OFFSET `DUALTIMER_OFFSET+16'h0024
`define DUALTIMER_TIMER2CONTROL_OFFSET `DUALTIMER_OFFSET+16'h0028
`define DUALTIMER_TIMER2INTCLR_OFFSET `DUALTIMER_OFFSET+16'h002C
`define DUALTIMER_TIMER2RIS_OFFSET `DUALTIMER_OFFSET+16'h0030
`define DUALTIMER_TIMER2MIS_OFFSET `DUALTIMER_OFFSET+16'h0034
`define DUALTIMER_TIMER2BGLOAD_OFFSET `DUALTIMER_OFFSET+16'h0038

`define APB_TEST_SLAVE_OFFSET 16'hB000
`define APB_TEST_SLAVE_DATA0_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0000
`define APB_TEST_SLAVE_DATA1_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0004
`define APB_TEST_SLAVE_DATA2_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0008
`define APB_TEST_SLAVE_DATA3_OFFSET `APB_TEST_SLAVE_OFFSET+16'h000C