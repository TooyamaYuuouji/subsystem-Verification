`ifndef AHBL_PKG_SV
`define AHBL_PKG_SV


`include "ahbl_interface.sv"

package ahbl_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "ahbl_defines.svh"
	`include "ahbl_types.sv"
	`include "ahbl_transaction.sv"
	`include "ahbl_agent_configuration.sv"
	`include "ahbl_mst_driver.sv"
	`include "ahbl_mst_monitor.sv"
	`include "ahbl_mst_sequencer.sv"
	`include "ahbl_mst_agent.sv"

endpackage : ahbl_pkg


`endif // AHBL_PKG_SV
