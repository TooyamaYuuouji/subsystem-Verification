
package ral_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "ral_timer.sv"

endpackage: ral_pkg
