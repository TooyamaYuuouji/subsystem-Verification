
package apb3_package;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "apb3_transaction.sv"
`include "apb3_configuration.sv"
`include "apb3_master_driver.sv"
`include "apb3_master_monitor.sv"
`include "apb3_master_sequencer.sv"
`include "apb3_master_agent.sv"

`include "apb3_master_base_seq.sv"

endpackage: apb3_package
