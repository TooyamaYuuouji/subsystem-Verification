`define TIMER0_OFFSET 16'h0000
`define TIMER0_CTRL_OFFSET `TIMER0_OFFSET+16'h0000
`define TIMER0_VALUE_OFFSET `TIMER0_OFFSET+16'h0004
`define TIMER0_RELOAD_OFFSET `TIMER0_OFFSET+16'h0008
`define TIMER0_INTCLEAR_OFFSET `TIMER0_OFFSET+16'h000C
`define TIMER0_IRQ 8

`define TIMER1_OFFSET 16'h1000
`define TIMER1_CTRL_OFFSET `TIMER1_OFFSET+16'h0000
`define TIMER1_VALUE_OFFSET `TIMER1_OFFSET+16'h0004
`define TIMER1_RELOAD_OFFSET `TIMER1_OFFSET+16'h0008
`define TIMER1_INTCLEAR_OFFSET `TIMER1_OFFSET+16'h000C
`define TIMER1_IRQ 9

`define DUALTIMER_OFFSET 16'h2000
`define DUALTIMER_TIMER1LOAD_OFFSET `DUALTIMER_OFFSET+16'h0000
`define DUALTIMER_TIMER1VALUE_OFFSET `DUALTIMER_OFFSET+16'h0004
`define DUALTIMER_TIMER1CONTROL_OFFSET `DUALTIMER_OFFSET+16'h0008
`define DUALTIMER_TIMER1INTCLR_OFFSET `DUALTIMER_OFFSET+16'h000C
`define DUALTIMER_TIMER1RIS_OFFSET `DUALTIMER_OFFSET+16'h0010
`define DUALTIMER_TIMER1MIS_OFFSET `DUALTIMER_OFFSET+16'h0014
`define DUALTIMER_TIMER1BGLOAD_OFFSET `DUALTIMER_OFFSET+16'h0018
`define DUALTIMER_TIMER2LOAD_OFFSET `DUALTIMER_OFFSET+16'h0020
`define DUALTIMER_TIMER2VALUE_OFFSET `DUALTIMER_OFFSET+16'h0024
`define DUALTIMER_TIMER2CONTROL_OFFSET `DUALTIMER_OFFSET+16'h0028
`define DUALTIMER_TIMER2INTCLR_OFFSET `DUALTIMER_OFFSET+16'h002C
`define DUALTIMER_TIMER2RIS_OFFSET `DUALTIMER_OFFSET+16'h0030
`define DUALTIMER_TIMER2MIS_OFFSET `DUALTIMER_OFFSET+16'h0034
`define DUALTIMER_TIMER2BGLOAD_OFFSET `DUALTIMER_OFFSET+16'h0038
`define DUALTIMER_IRQ 10

`define UART0_OFFSET 16'h4000
`define UART0_DATA_OFFSET `UART0_OFFSET+16'h0000
`define UART0_STATE_OFFSET `UART0_OFFSET+16'h0004
`define UART0_CTRL_OFFSET `UART0_OFFSET+16'h0008
`define UART0_INTCLEAR_OFFSET `UART0_OFFSET+16'h000C
`define UART0_BAUDDIV_OFFSET `UART0_OFFSET+16'h0010
`define UART0_RX_INT_IRQ 0
`define UART0_TX_INT_IRQ 1
`define UART0_OVERFLOW_INT_IRQ 12

`define UART1_OFFSET 16'h5000
`define UART1_DATA_OFFSET `UART1_OFFSET+16'h0000
`define UART1_STATE_OFFSET `UART1_OFFSET+16'h0004
`define UART1_CTRL_OFFSET `UART1_OFFSET+16'h0008
`define UART1_INTCLEAR_OFFSET `UART1_OFFSET+16'h000C
`define UART1_BAUDDIV_OFFSET `UART1_OFFSET+16'h0010
`define UART1_RX_INT_IRQ 2
`define UART1_TX_INT_IRQ 3
`define UART1_OVERFLOW_INT_IRQ 13

`define UART2_OFFSET 16'h6000
`define UART2_DATA_OFFSET `UART2_OFFSET+16'h0000
`define UART2_STATE_OFFSET `UART2_OFFSET+16'h0004
`define UART2_CTRL_OFFSET `UART2_OFFSET+16'h0008
`define UART2_INTCLEAR_OFFSET `UART2_OFFSET+16'h000C
`define UART2_BAUDDIV_OFFSET `UART2_OFFSET+16'h0010
`define UART2_RX_INT_IRQ 4
`define UART2_TX_INT_IRQ 5
`define UART2_OVERFLOW_INT_IRQ 14

`define APB_TEST_SLAVE_OFFSET 16'hB000
`define APB_TEST_SLAVE_DATA0_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0000
`define APB_TEST_SLAVE_DATA1_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0004
`define APB_TEST_SLAVE_DATA2_OFFSET `APB_TEST_SLAVE_OFFSET+16'h0008
`define APB_TEST_SLAVE_DATA3_OFFSET `APB_TEST_SLAVE_OFFSET+16'h000C