
package top_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import apb3_package::*;

`include "virtual_sequencer.sv"
// timer
`include "ral_timer.sv"
`include "timer_start_seq.sv"
`include "timer_clear_interrupt_seq.sv"
`include "timer_stop_seq.sv"

`include "scoreboard.sv"
`include "apb3_adapter.sv"
`include "base_env.sv"

`include "timer_base_test.sv"
`include "timer_test.sv"

endpackage: top_pkg
