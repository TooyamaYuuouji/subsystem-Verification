
package ral_pkg;

`include "ral_timer.sv"

endpackage: ral_pkg
